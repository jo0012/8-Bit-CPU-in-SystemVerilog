library verilog;
use verilog.vl_types.all;
entity bMux_tb is
end bMux_tb;
