library verilog;
use verilog.vl_types.all;
entity ControlUnit_tb is
end ControlUnit_tb;
