library verilog;
use verilog.vl_types.all;
entity Reg_8bit_tb is
end Reg_8bit_tb;
