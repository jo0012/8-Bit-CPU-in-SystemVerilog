library verilog;
use verilog.vl_types.all;
entity Top_level_tb is
end Top_level_tb;
