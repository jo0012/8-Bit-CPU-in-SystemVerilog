library verilog;
use verilog.vl_types.all;
entity PCnMUX_tb is
end PCnMUX_tb;
