library verilog;
use verilog.vl_types.all;
entity ROM_tb is
end ROM_tb;
